library IEEE;
use IEEE.STD_LOGIC_1164.all;



entity objects_draw is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   CLK  					: in std_logic;
		RESETn				: in std_logic;
		oCoord_X				: in integer;
		oCoord_Y				: in integer;
		bounce_type 		: out std_logic_vector(4 downto 0) ;
		drawing_request	: out std_logic ;
		mVGA_RGB 			: out std_logic_vector(7 downto 0) 
	);
end entity;

architecture behav of objects_draw is 

	constant no_bounce			 		: std_logic_vector (4 downto 0) := "00000";
	constant horizontal_floor 			: std_logic_vector (4 downto 0) := "00001";
	constant left_down_slope 			: std_logic_vector (4 downto 0) := "00010";
	constant left_vertical_wall 		: std_logic_vector (4 downto 0) := "00011";
	constant left_up_slope 				: std_logic_vector (4 downto 0) := "00100";
	constant horizontal_ceiling 		: std_logic_vector (4 downto 0) := "00101";
	constant right_up_slope 			: std_logic_vector (4 downto 0) := "00110";
	constant right_vertical_wall 		: std_logic_vector (4 downto 0) := "00111";
	constant right_down_slope 			: std_logic_vector (4 downto 0) := "01000";
	constant death				 		: std_logic_vector (4 downto 0) := "01001";

	--floor:
	constant floor_start_x 	: integer := 0;
	constant floor_start_y 	: integer := 450;
	constant floor_X_size 	: integer := 640;
	constant floor_Y_size 	: integer := 31;
	constant floor_color  	: std_logic_vector(7 downto 0) := x"13";
	constant floor_bounce_type : std_logic_vector(4 downto 0) := horizontal_floor;
	signal floor_end_x : integer;
	signal floor_end_y : integer;
	signal floor_drawing_X : std_logic := '0';
	signal floor_drawing_Y : std_logic := '0';
	signal floor_drawing_req : std_logic := '0';
	--/floor
	
	--right_wall:
	constant right_wall_start_x 	: integer := 610;
	constant right_wall_start_y 	: integer := 30;
	constant right_wall_X_size 	: integer := 31;
	constant right_wall_Y_size 	: integer := 420;
	constant right_wall_color  	: std_logic_vector(7 downto 0) := x"13";
	constant right_wall_bounce_type : std_logic_vector(4 downto 0) := right_vertical_wall;
	signal right_wall_end_x : integer;
	signal right_wall_end_y : integer;
	signal right_wall_drawing_X : std_logic := '0';
	signal right_wall_drawing_Y : std_logic := '0';
	signal right_wall_drawing_req : std_logic := '0';
	--/right_wall
	
	--left_wall:
	constant left_wall_start_x 	: integer := 0;
	constant left_wall_start_y 	: integer := 30;
	constant left_wall_X_size 	: integer := 31;
	constant left_wall_Y_size 	: integer := 420;
	constant left_wall_color  	: std_logic_vector(7 downto 0) := x"13";
	constant left_wall_bounce_type : std_logic_vector(4 downto 0) := left_vertical_wall;
	signal left_wall_end_x : integer;
	signal left_wall_end_y : integer;
	signal left_wall_drawing_X : std_logic := '0';
	signal left_wall_drawing_Y : std_logic := '0';
	signal left_wall_drawing_req : std_logic := '0';
	--/left_wall
	
	--ceiling:
	constant ceiling_start_x 	: integer := 0;
	constant ceiling_start_y 	: integer := 0;
	constant ceiling_X_size 	: integer := 640;
	constant ceiling_Y_size 	: integer := 31;
	constant ceiling_color  	: std_logic_vector(7 downto 0) := x"13";
	constant ceiling_bounce_type : std_logic_vector(4 downto 0) := horizontal_ceiling;
	signal ceiling_end_x : integer;
	signal ceiling_end_y : integer;
	signal ceiling_drawing_X : std_logic := '0';
	signal ceiling_drawing_Y : std_logic := '0';
	signal ceiling_drawing_req : std_logic := '0';
	--/ceiling
	
	--left_down_slope:
	constant left_down_slope_start_x 	: integer := 31;
	constant left_down_slope_start_y 	: integer := 282;
	constant left_down_slope_X_size 	: integer := 84;
	constant left_down_slope_Y_size 	: integer := 84;
	constant left_down_slope_color  	: std_logic_vector(7 downto 0) := x"13";
	constant left_down_slope_bounce_type : std_logic_vector(4 downto 0) := left_down_slope;
	signal left_down_slope_end_x : integer;
	signal left_down_slope_end_y : integer;
	signal left_down_slope_drawing_X : std_logic := '0';
	signal left_down_slope_drawing_Y : std_logic := '0';
	signal left_down_slope_drawing_req : std_logic := '0';
	signal left_down_slope_Coord_X : integer := 0;-- offset from start position 
	signal left_down_slope_Coord_Y : integer := 0;
	--/left_down_slope
	
	type left_down_slope_object_form is array (0 to left_down_slope_Y_size - 1 , 0 to left_down_slope_X_size - 1) of std_logic;
	constant left_down_slope_object : left_down_slope_object_form := (
("100000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("110000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111100000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111110000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111100000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111110000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111100000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111110000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111100000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111110000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111100000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111110000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111100000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111100000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111110000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111100000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111110000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111110000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111100000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111110000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111110000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111100000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111110000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111100000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111110000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111100000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111110000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111100000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111110000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111100000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111110000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111100000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111110000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111100000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111110000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111100000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111110000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111100000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111110000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111100000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111110000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111100000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111110000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111")

);
	
	--left_up_slope:
	constant left_up_slope_start_x 	: integer := 31;
	constant left_up_slope_start_y 	: integer := 31;
	constant left_up_slope_X_size 	: integer := 84;
	constant left_up_slope_Y_size 	: integer := 84;
	constant left_up_slope_color  	: std_logic_vector(7 downto 0) := x"13";
	constant left_up_slope_bounce_type : std_logic_vector(4 downto 0) := left_up_slope;
	signal left_up_slope_end_x : integer;
	signal left_up_slope_end_y : integer;
	signal left_up_slope_drawing_X : std_logic := '0';
	signal left_up_slope_drawing_Y : std_logic := '0';
	signal left_up_slope_drawing_req : std_logic := '0';
	signal left_up_slope_Coord_X : integer := 0;-- offset from start position 
	signal left_up_slope_Coord_Y : integer := 0;
	--/left_up_slope
	
	type left_up_slope_object_form is array (0 to left_up_slope_Y_size - 1 , 0 to left_up_slope_X_size - 1) of std_logic;
	constant left_up_slope_object : left_up_slope_object_form := (
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111110000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111100000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111110000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111100000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111110000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111100000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111110000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111100000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111110000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111100000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111110000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111100000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111110000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111100000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111110000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111100000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111110000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111100000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111110000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111100000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111110000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111100000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111110000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111110000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111100000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111110000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111110000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111100000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111110000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111100000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111100000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111110000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111101000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111110000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111100000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111110100000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111100000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111110000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111100000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111110000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111100000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("110000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);
	
	--right_down_slope:
	constant right_down_slope_start_x 	: integer := 365;
	constant right_down_slope_start_y 	: integer := 282;
	constant right_down_slope_X_size 	: integer := 84;
	constant right_down_slope_Y_size 	: integer := 84;
	constant right_down_slope_color  	: std_logic_vector(7 downto 0) := x"13";
	constant right_down_slope_bounce_type : std_logic_vector(4 downto 0) := right_down_slope;
	signal right_down_slope_end_x : integer;
	signal right_down_slope_end_y : integer;
	signal right_down_slope_drawing_X : std_logic := '0';
	signal right_down_slope_drawing_Y : std_logic := '0';
	signal right_down_slope_drawing_req : std_logic := '0';
	signal right_down_slope_Coord_X : integer := 0;-- offset from start position 
	signal right_down_slope_Coord_Y : integer := 0;
	--/right_down_slope
	
	type right_down_slope_object_form is array (0 to right_down_slope_Y_size - 1 , 0 to right_down_slope_X_size - 1) of std_logic;
	constant right_down_slope_object : right_down_slope_object_form := (
("000000000000000000000000000000000000000000000000000000000000000000000000000000000001"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000011"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000001111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000011111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000001111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000011111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000001111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000011111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000001111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000011111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000001111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000011111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000001111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000011111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000001111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000011111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000001111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000011111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000001111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000011111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000001111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000011111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000001111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000011111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000001111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000011111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000001111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000011111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000001111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000011111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000001111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000011111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000001111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000011111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000001111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000011111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000001111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000011111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000001111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000011111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000001111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000011111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000001111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000011111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000001111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000011111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000001111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000011111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000001111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000011111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000001111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000011111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111")
);

	
	--right_up_slope:
	constant right_up_slope_start_x 	: integer := 365;
	constant right_up_slope_start_y 	: integer := 31;
	constant right_up_slope_X_size 	: integer := 84;
	constant right_up_slope_Y_size 	: integer := 84;
	constant right_up_slope_color  	: std_logic_vector(7 downto 0) := x"13";
	constant right_up_slope_bounce_type : std_logic_vector(4 downto 0) := right_up_slope;
	signal right_up_slope_end_x : integer;
	signal right_up_slope_end_y : integer;
	signal right_up_slope_drawing_X : std_logic := '0';
	signal right_up_slope_drawing_Y : std_logic := '0';
	signal right_up_slope_drawing_req : std_logic := '0';
	signal right_up_slope_Coord_X : integer := 0;-- offset from start position 
	signal right_up_slope_Coord_Y : integer := 0;
	--/right_up_slope

	type right_up_slope_object_form is array (0 to right_up_slope_Y_size - 1 , 0 to right_up_slope_X_size - 1) of std_logic;
	constant right_up_slope_object : right_up_slope_object_form := (
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000011111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000001111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000011111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000001111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000011111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000001111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000011111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000001111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000011111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000001111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000011111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000001111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000011111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000001111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000011111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000001111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000011111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000001111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000011111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000001111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000011111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000001111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000011111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000001111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000011111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000001111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000011111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000001111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000011111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000001111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000011111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000001111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000011111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000001111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000011111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000001111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000011111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000001111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000011111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000001111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000011111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000001111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000011111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000001111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000011111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000001111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000011111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000001111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000011111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000001111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000011"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000001")
);	
	
	
	--right_middle_slope:
	constant right_middle_slope_start_x 	: integer := 449;
	constant right_middle_slope_start_y 	: integer := 115;
	constant right_middle_slope_X_size 	: integer := 84;
	constant right_middle_slope_Y_size 	: integer := 84;
	constant right_middle_slope_color  	: std_logic_vector(7 downto 0) := x"13";
	constant right_middle_slope_bounce_type : std_logic_vector(4 downto 0) := right_up_slope;
	signal right_middle_slope_end_x : integer;
	signal right_middle_slope_end_y : integer;
	signal right_middle_slope_drawing_X : std_logic := '0';
	signal right_middle_slope_drawing_Y : std_logic := '0';
	signal right_middle_slope_drawing_req : std_logic := '0';
	signal right_middle_slope_Coord_X : integer := 0;-- offset from start position 
	signal right_middle_slope_Coord_Y : integer := 0;
	--/right_up_slope
	
	type right_middle_slope_object_form is array (0 to right_middle_slope_Y_size - 1 , 0 to right_middle_slope_X_size - 1) of std_logic;
	constant right_middle_slope_object : right_middle_slope_object_form := (
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000011111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000001111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000011111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000001111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000011111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000001111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000011111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000001111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000011111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000001111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000011111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000001111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000011111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000001111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000011111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000001111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000011111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000001111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000011111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000001111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000011111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000001111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000011111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000001111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000011111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000001111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000011111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000001111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000011111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000001111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000011111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000001111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000011111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000001111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000011111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000001111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000011111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000001111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000011111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000001111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000011111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000001111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000011111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000001111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000011111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000001111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000011111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000001111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000011111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000001111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000011"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000001")
);	



--stage_left:
	constant stage_left_start_x 	: integer := 0;
	constant stage_left_start_y 	: integer := 450;
	constant stage_left_X_size 	: integer := 640;
	constant stage_left_Y_size 	: integer := 31;
	constant stage_left_color  	: std_logic_vector(7 downto 0) := x"13";
	constant stage_left_bounce_type : std_logic_vector(4 downto 0) := horizontal_floor;
	signal stage_left_end_x : integer;
	signal stage_left_end_y : integer;
	signal stage_left_drawing_X : std_logic := '0';
	signal stage_left_drawing_Y : std_logic := '0';
	signal stage_left_drawing_req : std_logic := '0';
--/stage_left

--stage_right:
	constant stage_right_start_x 	: integer := 0;
	constant stage_right_start_y 	: integer := 450;
	constant stage_right_X_size 	: integer := 640;
	constant stage_right_Y_size 	: integer := 31;
	constant stage_right_color  	: std_logic_vector(7 downto 0) := x"13";
	constant stage_right_bounce_type : std_logic_vector(4 downto 0) := horizontal_floor;
	signal stage_right_end_x : integer;
	signal stage_right_end_y : integer;
	signal stage_right_drawing_X : std_logic := '0';
	signal stage_right_drawing_Y : std_logic := '0';
	signal stage_right_drawing_req : std_logic := '0';
--/stage_right

--tunnel_wall:
	constant tunnel_wall_start_x 	: integer := 0;
	constant tunnel_wall_start_y 	: integer := 450;
	constant tunnel_wall_X_size 	: integer := 640;
	constant tunnel_wall_Y_size 	: integer := 31;
	constant tunnel_wall_color  	: std_logic_vector(7 downto 0) := x"13";
	constant tunnel_wall_bounce_type : std_logic_vector(4 downto 0) := horizontal_floor;
	signal tunnel_wall_end_x : integer;
	signal tunnel_wall_end_y : integer;
	signal tunnel_wall_drawing_X : std_logic := '0';
	signal tunnel_wall_drawing_Y : std_logic := '0';
	signal tunnel_wall_drawing_req : std_logic := '0';
--/tunnel_wall
	
	
	--All Purpose :
	signal sig_draw_req : std_logic := '0';
	signal sig_draw_data: std_logic_vector (7 downto 0);
	signal sig_bounce_type : std_logic_vector (4 downto 0);
	--signal bCoord_X : integer := 0;-- offset from start position 
	--signal bCoord_Y : integer := 0;

	

--		


begin

	-- Calculate objects end boundaries
	left_down_slope_end_x	<= left_down_slope_X_size + left_down_slope_start_x;
	left_down_slope_end_y	<= left_down_slope_Y_size + left_down_slope_start_y;
	
	left_up_slope_end_x	<= left_up_slope_X_size + left_up_slope_start_x;
	left_up_slope_end_y	<= left_up_slope_Y_size + left_up_slope_start_y;
	
	right_down_slope_end_x	<= right_down_slope_X_size + right_down_slope_start_x;
	right_down_slope_end_y	<= right_down_slope_Y_size + right_down_slope_start_y;
	
	right_up_slope_end_x	<= right_up_slope_X_size + right_up_slope_start_x;
	right_up_slope_end_y	<= right_up_slope_Y_size + right_up_slope_start_y;
	
	right_middle_slope_end_x	<= right_middle_slope_X_size + right_middle_slope_start_x;
	right_middle_slope_end_y	<= right_middle_slope_Y_size + right_middle_slope_start_y;
	---------------------------------------------------------------
	
	
	floor_end_x	<= floor_X_size + floor_start_x;
	floor_end_y	<= floor_Y_size + floor_start_y;
	
	ceiling_end_x	<= ceiling_X_size + ceiling_start_x;
	ceiling_end_y	<= ceiling_Y_size + ceiling_start_y;
	
	left_wall_end_x	<= left_wall_X_size + left_wall_start_x;
	left_wall_end_y	<= left_wall_Y_size + left_wall_start_y;
	
	right_wall_end_x	<= right_wall_X_size + right_wall_start_x;
	right_wall_end_y	<= right_wall_Y_size + right_wall_start_y;
	
	------------------------------------------------------------------
	
	
	-- test if ooCoord is in the rectangle defined by Start and End 
	floor_drawing_X	<= '1' when  (oCoord_X  >= floor_start_x) and  (oCoord_X < floor_end_x) else '0';
   floor_drawing_Y	<= '1' when  (oCoord_Y  >= floor_start_y) and  (oCoord_Y < floor_end_y) else '0';
	
	ceiling_drawing_X	<= '1' when  (oCoord_X  >= ceiling_start_x) and  (oCoord_X < ceiling_end_x) else '0';
   ceiling_drawing_Y	<= '1' when  (oCoord_Y  >= ceiling_start_y) and  (oCoord_Y < ceiling_end_y) else '0';
	
	left_wall_drawing_X	<= '1' when  (oCoord_X  >= left_wall_start_x) and  (oCoord_X < left_wall_end_x) else '0';
   left_wall_drawing_Y	<= '1' when  (oCoord_Y  >= left_wall_start_y) and  (oCoord_Y < left_wall_end_y) else '0';
	
	right_wall_drawing_X	<= '1' when  (oCoord_X  >= right_wall_start_x) and  (oCoord_X < right_wall_end_x) else '0';
   right_wall_drawing_Y	<= '1' when  (oCoord_Y  >= right_wall_start_y) and  (oCoord_Y < right_wall_end_y) else '0';	
	--------------------------------------------------------------------------------------------------------
	
   	left_down_slope_drawing_X	<= '1' when  (oCoord_X  >= left_down_slope_start_x) and  (oCoord_X < left_down_slope_end_x) else '0';
   left_down_slope_drawing_Y	<= '1' when  (oCoord_Y  >= left_down_slope_start_y) and  (oCoord_Y < left_down_slope_end_y) else '0';
	
   	left_up_slope_drawing_X	<= '1' when  (oCoord_X  >= left_up_slope_start_x) and  (oCoord_X < left_up_slope_end_x) else '0';
   left_up_slope_drawing_Y	<= '1' when  (oCoord_Y  >= left_up_slope_start_y) and  (oCoord_Y < left_up_slope_end_y) else '0';
	
   	right_down_slope_drawing_X	<= '1' when  (oCoord_X  >= right_down_slope_start_x) and  (oCoord_X < right_down_slope_end_x) else '0';
   right_down_slope_drawing_Y	<= '1' when  (oCoord_Y  >= right_down_slope_start_y) and  (oCoord_Y < right_down_slope_end_y) else '0';
	
   	right_up_slope_drawing_X	<= '1' when  (oCoord_X  >= right_up_slope_start_x) and  (oCoord_X < right_up_slope_end_x) else '0';
   right_up_slope_drawing_Y	<= '1' when  (oCoord_Y  >= right_up_slope_start_y) and  (oCoord_Y < right_up_slope_end_y) else '0';

-- calculate offset from start corner 
	left_down_slope_Coord_X 	<= (oCoord_X - left_down_slope_start_x) when ( left_down_slope_drawing_X = '1' and  left_down_slope_drawing_Y = '1'  ) else 0 ; 
	left_down_slope_Coord_Y 	<= (oCoord_Y - left_down_slope_start_y) when ( left_down_slope_drawing_X = '1' and  left_down_slope_drawing_Y = '1'  ) else 0 ;
	
	left_up_slope_Coord_X 	<= (oCoord_X - left_up_slope_start_x) when ( left_up_slope_drawing_X = '1' and  left_up_slope_drawing_Y = '1'  ) else 0 ; 
	left_up_slope_Coord_Y 	<= (oCoord_Y - left_up_slope_start_y) when ( left_up_slope_drawing_X = '1' and  left_up_slope_drawing_Y = '1'  ) else 0 ;
	
	right_down_slope_Coord_X 	<= (oCoord_X - right_down_slope_start_x) when ( right_down_slope_drawing_X = '1' and  right_down_slope_drawing_Y = '1'  ) else 0 ; 
	right_down_slope_Coord_Y 	<= (oCoord_Y - right_down_slope_start_y) when ( right_down_slope_drawing_X = '1' and  right_down_slope_drawing_Y = '1'  ) else 0 ;
	
	right_up_slope_Coord_X 	<= (oCoord_X - right_up_slope_start_x) when ( right_up_slope_drawing_X = '1' and  right_up_slope_drawing_Y = '1'  ) else 0 ; 
	right_up_slope_Coord_Y 	<= (oCoord_Y - right_up_slope_start_y) when ( right_up_slope_drawing_X = '1' and  right_up_slope_drawing_Y = '1'  ) else 0 ;

	right_middle_slope_Coord_X 	<= (oCoord_X - right_middle_slope_start_x) when ( right_middle_slope_drawing_X = '1' and  right_middle_slope_drawing_Y = '1'  ) else 0 ; 
	right_middle_slope_Coord_Y 	<= (oCoord_Y - right_middle_slope_start_y) when ( right_middle_slope_drawing_X = '1' and  right_middle_slope_drawing_Y = '1'  ) else 0 ;

	
process ( RESETn, CLK)

  		
   begin
	
	
	
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

	elsif rising_edge(CLK) then
	
		sig_draw_req <= '0';
		sig_bounce_type <= no_bounce;
		if ( (floor_drawing_X ='1') and (floor_drawing_Y = '1') ) then
			sig_draw_req <= '1';
			sig_draw_data <= floor_color;
			sig_bounce_type <= floor_bounce_type;
		end if;
		

		if ((ceiling_drawing_X ='1') and (ceiling_drawing_Y = '1') ) then
			sig_draw_req <= '1';
			sig_draw_data <= ceiling_color;
			sig_bounce_type <= ceiling_bounce_type;
		end if;	
		

		if ((left_wall_drawing_X ='1') and (left_wall_drawing_Y = '1')) then
			sig_draw_req <= '1';
			sig_draw_data <= left_wall_color;
			sig_bounce_type <= left_wall_bounce_type;
		end if;

		if ((right_wall_drawing_X ='1') and (right_wall_drawing_Y = '1')) then
			sig_draw_req <= '1';
			sig_draw_data <= right_wall_color;
			sig_bounce_type <= right_wall_bounce_type;
		end if;
		
		----------------------------------------------------------------------------
		
		if ((left_down_slope_drawing_X ='1') and (left_down_slope_drawing_Y = '1')) then
			sig_draw_req <= left_down_slope_object(left_down_slope_Coord_Y,left_down_slope_Coord_X);
			sig_draw_data <= left_down_slope_color;
			if left_down_slope_object(left_down_slope_Coord_Y,left_down_slope_Coord_X) = '1' then
				sig_bounce_type <= left_down_slope_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;
		
		if ((left_up_slope_drawing_X ='1') and (left_up_slope_drawing_Y = '1')) then
			sig_draw_req <= left_up_slope_object(left_up_slope_Coord_Y,left_up_slope_Coord_X);
			sig_draw_data <= left_up_slope_color;
			if left_up_slope_object(left_up_slope_Coord_Y,left_up_slope_Coord_X) = '1' then
				sig_bounce_type <= left_up_slope_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;
		
		if ((right_down_slope_drawing_X ='1') and (right_down_slope_drawing_Y = '1')) then
			sig_draw_req <= right_down_slope_object(right_down_slope_Coord_Y, right_down_slope_Coord_X);
			sig_draw_data <= right_down_slope_color;
			if right_down_slope_object(right_down_slope_Coord_Y, right_down_slope_Coord_X) = '1' then
				sig_bounce_type <= right_down_slope_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;
		
		if ((right_up_slope_drawing_X ='1') and (right_up_slope_drawing_Y = '1')) then
			sig_draw_req <= right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_Coord_X);
			sig_draw_data <= right_up_slope_color;
			if right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_Coord_X) = '1' then
				sig_bounce_type <= right_up_slope_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;
		
		if ((right_middle_slope_drawing_X ='1') and (right_middle_slope_drawing_Y = '1')) then
			sig_draw_req <= right_middle_slope_object(right_middle_slope_Coord_Y,right_middle_slope_Coord_X);
			sig_draw_data <= right_middle_slope_color;
			if right_middle_slope_object(right_middle_slope_Coord_Y,right_middle_slope_Coord_X) = '1' then
				sig_bounce_type <= right_middle_slope_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		----------------------------------------------------------------------------
	
			mVGA_RGB	<=  sig_draw_data;	--get from colors table 
			drawing_request	<=  sig_draw_req ; -- get from mask table if inside rectangle
			bounce_type <= sig_bounce_type;
	end if;

  end process;

		
end architecture;	